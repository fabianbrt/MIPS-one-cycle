----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/12/2025 09:21:48 PM
-- Design Name: 
-- Module Name: SSD_pali - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SSD_pali is
    Port ( digits : in STD_LOGIC_VECTOR (31 downto 0);
       clk : in STD_LOGIC;
       cat : out STD_LOGIC_VECTOR (6 downto 0);
       an : out STD_LOGIC_VECTOR (7 downto 0));
end SSD_pali;

architecture Behavioral of SSD_pali is

begin


end Behavioral;
